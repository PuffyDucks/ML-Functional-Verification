module mod (
    input [7:0] a,
    output [5:0] result
);

    assign result = a[5:0];

endmodule
